module regfile(input clk, rst, we3,
               input  [4:0]  ra1, ra2, wa3, 
               input  [31:0] wd3, 
               output [31:0] rd1, rd2);

  	reg [31:0] rf [31:0];

	always@(posedge rst) begin
		rf[0] <= 32'h00000000;
		rf[1] <= 32'h00000000;
		rf[2] <= 32'h00000000;
		rf[3] <= 32'h00000000;
		rf[4] <= 32'h00000000;
		rf[5] <= 32'h00000000;
		rf[6] <= 32'h00000000;
		rf[7] <= 32'h00000000;
		rf[8] <= 32'h00000000;						
		rf[9] <= 32'h00000000;						
		rf[10] <= 32'h00000000;
		rf[11] <= 32'h00000000;
		rf[12] <= 32'h00000000;
		rf[13] <= 32'h00000000;
		rf[14] <= 32'h00000000;
		rf[15] <= 32'h00000000;
		rf[16] <= 32'h00000000;
		rf[17] <= 32'h00000000;
		rf[18] <= 32'h00000000;					
		rf[19] <= 32'h00000000;					
		rf[20] <= 32'h00000000;					
		rf[21] <= 32'h00000000;
		rf[22] <= 32'h00000000;					
		rf[23] <= 32'h00000000;
		rf[24] <= 32'h00000000;
		rf[25] <= 32'h00000000;
		rf[26] <= 32'h00000000;
		rf[27] <= 32'h00000000;
		rf[28] <= 32'h00000000;
		rf[29] <= 32'h00000000;
		rf[30] <= 32'h00000000;
		rf[31] <= 32'h00000000;
	end

  	always @(negedge clk) begin
   		if (we3 & rst == 0) begin
			rf[wa3] <= wd3;	
		end
	end
  	assign rd1 = (ra1 != 0) ? rf[ra1] : 0;
  	assign rd2 = (ra2 != 0) ? rf[ra2] : 0;
endmodule